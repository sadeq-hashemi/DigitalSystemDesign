module barcode(clk, rst_n, BC, clr_ID_vld, ID, ID_vld); 

input clk, rst_n
input BC, clr_ID_vld; 
output [7:0] ID; 
output ID_vld; 

reg  
reg 
localparam byte_done 4'b1000



endmodule
